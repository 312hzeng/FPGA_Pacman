module food(input Reset, input clock,
				input [9:0] PacmanX, PacmanY, DrawX, DrawY,
			   output isFood, finish);
	logic food[29][28];
	
	int food_array[812];
	logic [5:0] pacmanx, pacmany, drawx, drawy;
	assign food_array ='{ 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //0
								 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //1
								 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, ///0
								 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //3
								 0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,0, //4
								 0,0,1,0,0,0,1,0,0,0,0,0,1,1,0,1,0,0,0,0,0,0,1,0,0,0,1,0, //5
								 0,0,1,0,0,0,1,0,0,0,0,0,1,1,0,1,0,0,0,0,0,0,1,0,0,0,1,0, //6
								 0,0,1,0,0,0,1,0,0,0,0,0,1,1,0,1,0,0,0,0,0,0,1,0,0,0,1,0, //7
								 0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0, //8
								 0,0,1,0,0,0,1,0,1,1,1,0,0,0,0,0,0,0,1,1,1,0,1,0,0,0,1,0, //9
								 0,0,1,1,1,1,1,0,1,1,1,1,1,1,0,1,1,1,1,1,1,0,1,1,1,1,1,0, //01
								 0,0,0,0,0,0,1,0,0,0,0,0,1,1,0,1,1,0,0,0,0,0,1,0,0,0,0,0, //00
								 0,0,0,0,0,0,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,0,0,0,0,0, //00
								 0,0,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,0, //03 
								 0,0,0,0,0,0,1,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,1,0,0,0,0,0, //04
								 0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0, //05
								 0,0,0,0,0,0,1,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,1,0,0,0,0,0, //06
								 0,0,0,0,0,0,1,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,1,0,0,0,0,0, //07
								 0,0,1,1,1,1,1,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,1,1,1,1,1,0, //08
								 0,0,0,0,0,0,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,0,0,0,0,0, //09
								 0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0, //01
								 0,0,1,0,0,0,1,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,1,0,0,0,1,0, //00
								 0,0,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,0, //00
								 0,0,1,1,1,0,1,1,0,1,0,0,0,0,0,0,0,0,0,1,0,1,1,0,1,1,1,0, //03
								 0,0,0,0,1,0,1,1,0,1,1,1,1,1,0,1,1,1,1,1,0,1,1,0,1,0,0,0, //04
								 0,0,1,1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1,1,0, //05
								 0,0,1,1,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,1,1,0, //06
								 0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0, //07 
								 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0 
								 };  //08
													
				
	always_ff @ (posedge Reset or posedge clock )
   begin
		if(Reset)
		begin
			for(int i = 0; i < 29; i++)
			begin
				for(int j = 0; j < 28; j++)
				begin
					food[i][j] <= food_array[i * 28 + j];
				end
			end
		end
		
		
		else
		begin
			 pacmanx = PacmanX[9:4];
			 pacmany = PacmanY[9:4];
		    if(pacmanx <= 27 && pacmanx >= 0 && pacmany <= 28 && pacmany >= 0)
				food[pacmany][pacmanx] <= 0;
		end
	
	end

	always_comb
	begin
	drawx = DrawX[9:4];
	drawy = DrawY[9:4];
	if(drawx <= 27 && drawx >= 0 && drawy <= 28 && drawy >= 0 && food[drawy][drawx] == 1 )
	begin
			isFood = 1'b1;
	end
	else
			isFood = 1'b0;
	end
	
	always_comb
	begin
		finish = 1;
		for(int i = 0; i < 29; i++)
			begin
				for(int j = 0; j < 28; j++)
				begin
					if(food[i][j] == 1)
						finish = 0;
				end
			end
	end
endmodule
