module intro (input [9:0]DrawX,
             input [9:0] DrawY,
             output [1:0]intro
				 );
								  
	 
	 
	 always_comb 
	 begin
	    logic [10:0]index;
		 logic [5:0] drawx, drawy;
		 
		 int maze[900]; //30 * 30
		 maze = '{
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //0
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //1
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //2
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //3
			 0,1,1,1,1,2,2,2,2,3,3,3,3,0,0,0,1,0,0,0,1,2,2,2,2,3,0,0,3,0, //4
			 0,1,0,0,1,2,0,0,2,3,0,0,0,0,0,0,1,1,0,1,1,2,0,0,2,3,3,0,3,0, //5
			 0,1,0,0,1,2,0,0,2,3,0,0,0,0,0,0,1,1,1,1,1,2,0,0,2,3,3,0,3,0, //6
			 0,1,1,1,1,2,0,0,2,3,0,0,0,0,0,0,1,0,1,0,1,2,0,0,2,3,3,0,3,0, //7
			 0,1,0,0,0,2,0,0,2,3,0,0,0,0,0,0,1,0,1,0,1,2,0,0,2,3,3,0,3,0, //8
			 0,1,0,0,0,2,2,2,2,3,0,0,0,1,1,0,1,0,0,0,1,2,2,2,2,3,0,3,3,0, //9
			 0,1,0,0,0,2,0,0,2,3,0,0,0,0,0,0,1,0,0,0,1,2,0,0,2,3,0,3,3,0, //10
			 0,1,0,0,0,2,0,0,2,3,0,0,0,0,0,0,1,0,0,0,1,2,0,0,2,3,0,3,3,0, //11
			 0,1,0,0,0,2,0,0,2,3,0,0,0,0,0,0,1,0,0,0,1,2,0,0,2,3,0,3,3,0, //12
			 0,1,0,0,0,2,0,0,2,3,3,3,3,0,0,0,1,0,0,0,1,2,0,0,2,3,0,0,3,0, //13 
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //14
			 0,1,1,1,2,2,2,3,3,3,2,2,2,1,1,1,0,0,1,0,1,2,2,2,3,0,3,0,1,0, //15
			 0,1,0,1,2,0,2,3,0,0,2,0,0,1,0,0,0,0,1,1,0,2,0,0,3,3,3,1,1,0, //16
			 0,1,1,1,2,2,2,3,3,3,2,2,2,1,1,1,0,0,1,1,0,2,2,2,0,3,0,0,1,0, //17
			 0,1,0,0,2,2,0,3,0,0,0,0,2,0,0,1,0,0,1,1,0,2,0,0,0,3,0,0,1,0, //18
			 0,1,0,0,2,0,2,3,3,3,2,2,2,1,1,1,0,0,1,0,1,2,2,2,0,3,0,1,1,1, //19
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //20
			 0,1,1,1,2,2,2,0,0,3,3,3,1,1,1,2,2,2,1,1,1,2,2,2,0,0,3,3,0,0, //21
			 0,0,1,0,2,0,2,0,0,3,0,0,0,1,0,2,0,2,1,0,1,0,2,0,0,0,3,3,0,0, //22
			 0,0,1,0,2,0,2,0,0,3,3,3,0,1,0,2,2,2,1,1,1,0,2,0,0,0,3,3,0,0, //23
			 0,0,1,0,2,0,2,0,0,0,0,3,0,1,0,2,0,2,1,1,0,0,2,0,0,0,0,0,0,0, //24
			 0,0,1,0,2,2,2,0,0,3,3,3,0,1,0,2,0,2,1,0,1,0,2,0,0,0,3,3,0,0, //25
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //26
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //27 
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, //28
			 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0 //29
		 };
	
	    drawx[5:0] = DrawX[9:4];
		 drawy[5:0] = DrawY[9:4];

	 if(drawx <= 29 && drawx >= 0 && drawy <= 29 && drawy >= 0)
		 begin
	        index = drawy * 30 + drawx;
			  if(maze[index] == 1)
			      intro = 1;
			  else if(maze[index] == 2)
						intro = 2;
			  else if(maze[index] == 3)
						intro = 3;
			  else
					intro = 0;
		 end
		 
		 else
		     intro = 0;
	 end
endmodule
